`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// Engineer: 		 Balazs Nagy
// 
// Create Date:    01:02:49 06/19/2015 
// Module Name:    draw_strings  
// Project Name: 	 Tetris Game
// Description:	 Draw Strings for the Tetris game
//	
//////////////////////////////////////////////////////////////////////////////////
module draw_strings(
    input vga_clk,
    input rst,
    input [10:0] x,
    input [9:0] y,
    output [1:0] r,
    output [1:0] g,
    output [1:0] b,
    output reg dav
);



endmodule
